module MainModule();


endmodule
