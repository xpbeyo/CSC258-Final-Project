module MainModule(dir);
    input [1:0] dir;

endmodule
